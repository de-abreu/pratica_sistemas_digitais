library ieee;
use ieee.std_logic_1164.all;

package array_t is
    type vector_array is array (natural range <>) of STD_LOGIC_VECTOR;
end package array_t;
