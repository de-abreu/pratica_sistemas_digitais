library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.state_t.all;

entity testbench is
end testbench;

architecture Behavioral of testbench is

    -- Component declaration for the segment_counter
    component segment_counter_one_hot is
    port (
        input, clk, rst : in  std_logic := '0';
        output          : out std_logic;
        s               : out state
     );
    end component;

    -- Signals for the testbench
    signal input, clk, rst, output  : std_logic := '0';
    signal s : state;

    -- Clock period constant
    constant clk_period : time := 10 ns;

begin

    -- Instantiate the segment_counter unit under test (UUT)
    uut : segment_counter_one_hot
    port map (
        input => input,
        clk => clk,
        rst => rst,
        output => output,
        s => s
    );

    -- Clock generation process
    clk_process : process
    begin
        wait for clk_period / 2;
        clk <= not clk;
    end process;

    -- Test process to simulate different conditions
    test_process : process
    begin
        -- Initial reset
        rst <= '0';
        wait for clk_period * 2;
        rst <= '1';
        wait for clk_period * 2;

        -- Test 1: Segment shorter than 4 bits (3 bits of '0')
        input <= '0';
        wait for clk_period * 3;  -- 3 cycles of '0'
        input <= '1';  -- Change to break the segment
        assert output = '0' report "Failed: Output should be '0' for segment < 4 bits (0s)" severity error;
        wait for clk_period * 2;

        -- Test 2: Segment shorter than 4 bits (3 bits of '1')
        input <= '1';
        wait for clk_period * 3;  -- 3 cycles of '1'
        input <= '0';  -- Change to break the segment
        assert output = '0' report "Failed: Output should be '0' for segment < 4 bits (1s)" severity error;
        wait for clk_period * 2;

        -- Test 3: Segment exactly 4 bits (4 bits of '0')
        input <= '0';
        wait for clk_period * 4;  -- 4 cycles of '0'
        assert output = '1' report "Failed: Output should be '1' for segment = 4 bits (0s)" severity error;
        wait for clk_period * 2;

        -- Test 4: Segment exactly 4 bits (4 bits of '1')
        input <= '1';
        wait for clk_period * 4;  -- 4 cycles of '1'
        assert output = '1' report "Failed: Output should be '1' for segment = 4 bits (1s)" severity error;
        wait for clk_period * 2;

        -- Test 5: Reset test
        rst <= '0';
        wait for clk_period * 2;
        assert output = '0' report "Failed: Output should be '0' after reset" severity error;
        rst <= '1';
        wait for clk_period * 2;

        -- End of simulation
        report "All tests completed successfully" severity note;
        wait;
    end process;

end Behavioral;
