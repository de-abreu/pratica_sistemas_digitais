library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.arrays_t.all;
use work.instructions_t.all;

entity cpu_tb is
end entity cpu_tb;

architecture Behaviour of cpu_tb is
    -- CPU signams
begin
end rchitecture Behaviour
